module bcd7seg(
    input [3:0] b,
    output reg [7:0] h
);

//    _7_
//  2|   |6
//   |_1_|
//  3|   |5 
//   |_4_|.0

always@(*)
    case(b)
        4'd0:    h = ~(8'b11111101);//0  
        4'd1:    h = ~(8'b01100001);//1
        4'd2:    h = ~(8'b11011011);//2
        4'd3:    h = ~(8'b11110011);//3
        4'd4:    h = ~(8'b01100111);//4
        4'd5:    h = ~(8'b10110111);//5
        4'd6:    h = ~(8'b10111111);//6
        4'd7:    h = ~(8'b11100001);//7
        4'd8:    h = ~(8'b11111111);//8
        4'd9:    h = ~(8'b11110111);//9
        4'd10:   h = ~(8'b11101111);//A
        4'd11:   h = ~(8'b00111111);//b
        4'd12:   h = ~(8'b10011101);//C
        4'd13:   h = ~(8'b01111011);//d
        4'd14:   h = ~(8'b00111111);//E
        4'd15:   h = ~(8'b10001111);//F
        default: h = ~(8'b11111111);//8.
    endcase

endmodule



