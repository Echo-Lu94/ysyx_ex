module bcd7seg(
    input [4:0] b,
    output reg [7:0] h
);

//    _7_
//  2|   |6
//   |_1_|
//  3|   |5 
//   |_4_|.0

always@(*)
    case(b)
        5'd0:    h = ~(8'b11111100);//0  
        5'd1:    h = ~(8'b01100000);//1
        5'd2:    h = ~(8'b11011010);//2
        5'd3:    h = ~(8'b11110010);//3
        5'd4:    h = ~(8'b01100110);//4
        5'd5:    h = ~(8'b10110110);//5
        5'd6:    h = ~(8'b10111110);//6
        5'd7:    h = ~(8'b11100000);//7
        5'd8:    h = ~(8'b11111110);//8
        5'd9:    h = ~(8'b11110110);//9
        5'd10:   h = ~(8'b11101110);//A
        5'd11:   h = ~(8'b00111110);//b
        5'd12:   h = ~(8'b10011100);//C
        5'd13:   h = ~(8'b01111010);//d
        5'd14:   h = ~(8'b10011110);//E
        5'd15:   h = ~(8'b10001110);//F
//        default: h = ~(8'b11111110);//8.
        default: h = ~(8'b00000000);//light off
    endcase

endmodule



